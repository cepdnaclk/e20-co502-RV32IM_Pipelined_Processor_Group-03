module instruction_memory(
    input CLK,
    in 
);