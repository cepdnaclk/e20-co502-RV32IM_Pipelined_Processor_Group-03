module instruction_memory(
    input  clk,
    input [31:0] PC,
    input reset,

    output reg [31:0] instruction
);
    reg [31:0] memory [0:1023];
    integer i;

    // initial begin
    //     memory[0] = 32'b00000000001000001_000_00011_0110011; //ADD x3, x1, x2
    //     memory[1] = 32'b0100000_00010_00001_000_00100_0110011; //SUB x2, x1, x2
    //     memory[2] = 32'b00000000001100000010000000100011; //SW x3, 6(x0)
    //     memory[3] = 32'b00000000010000000010001000100011; //SW x4, 4(x0)
    //     memory[4] = 32'b00000000000000000010001010000011; //LW x2, 0(x0)
    //     memory[5] = 32'b00000000010000000010001100000011; //LW x1, 4(x0)
    //     memory[6] = 32'b000000001010_00100_000_00001_0010011; //ADDI x1, x4, 10
    //     memory[7] = 32'b000000000101_00100_000_00010_0010011; //ADDI x2, x4, 5
    // end

    //Instructions to check load use hazards    
    initial begin
        memory[0] = 32'b0000000_00010_00001_000_00011_0110011; //ADD x3, x1, x2
        memory[1] = 32'b0000000_00011_00001_000_00100_0110011; //ADD x4, x1, x3
    end

    //Fibb  0, 1, 1, 2, 3, 5, 8, 13
    // initial begin
    //     memory[0] = 32'b00000000000100000000000000010011;
    //     memory[1] = 32'b00000000000100001000000010010011; 
    //     memory[2] = 32'b00000000000000101000001010010011; 
    //     memory[3] = 32'b00000000000100000000000100110011; 
    //     memory[4] = 32'b00000000000000001000000000010011;
    //     memory[5] = 32'b00000000000000010000000010010011; 
    //     memory[6] = 32'b00000000001000000010001010100011; 
    //     memory[7] = 32'b00000000000000000000000000000000;
    //     memory[8] = 32'b00000000000000000000000000000000;
    //     memory[9] = 32'b00000000000000000000000000000000; 
    //     memory[10] = 32'b00000000010100000010001100000011;
    //     memory[11] = 32'b11111101110111111111001011101111; 

    // end

    always @(posedge clk) begin
        instruction <= memory[PC/4];
    end
endmodule