module register_file(data1,data2,addr1,addr2,write_enable,clk,reg_write_data,reset,write_reg_addr);
    input [4:0] addr1,addr2,write_reg_addr;
    input [31:0] reg_write_data;
    input R,clk,reset,write_enable;
    output [31:0] data1,data2;

    reg [31:0] register [31:0];

    assign data1 = register[addr1];
    assign data2 = register[addr2];

    always @ (posedge clk)
    begin
      if (reset == 1)
        begin
        register[0] <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        register[1] <= 32'b0000_0000_0000_0000_0000_0000_0000_0111;
        register[2] <= 32'b0000_0000_0000_0000_0000_0000_0000_0010;
        register[3] <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        register[4] <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        register[5] <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        register[6] <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        register[7] <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        register[8] <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        register[9] <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        register[10] <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        register[11] <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        register[12] <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        register[13] <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        register[14] <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        register[15] <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        register[16] <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        register[17] <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        register[18] <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        register[19] <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        register[20] <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        register[21] <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        register[22] <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        register[23] <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        register[24] <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        register[25] <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        register[26] <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        register[27] <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        register[28] <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        register[29] <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        register[30] <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        register[31] <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
        end
      else
        begin
          if (write_enable == 1)
            begin
                register[write_reg_addr] <= reg_write_data;
            end
        end
    end
endmodule